module processor (
    
);
    
endmodule
